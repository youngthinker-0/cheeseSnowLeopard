`include "lib/defines.vh"
module IF(
    input wire clk,
    input wire rst,
    input wire [`StallBus-1:0] stall,

    // input wire flush,
    // input wire [31:0] new_pc,

    input wire [`BR_WD-1:0] br_bus, // BR zongxian

    output wire [`IF_TO_ID_WD-1:0] if_to_id_bus, 

    output wire inst_sram_en,
    output wire [3:0] inst_sram_wen,
    output wire [31:0] inst_sram_addr,
    output wire [31:0] inst_sram_wdata
);
    reg [31:0] pc_reg;
    reg ce_reg;
    wire [31:0] next_pc;
    wire br_e;
    wire [31:0] br_addr;

    assign {
        br_e,
        br_addr 
    } = br_bus;


    always @ (posedge clk) begin
        if (rst) begin // start
            pc_reg <= 32'hbfbf_fffc;
        end
        else if (stall[0]==`NoStop) begin //next pc
            pc_reg <= next_pc;
        end
    end

    always @ (posedge clk) begin
        if (rst) begin //
            ce_reg <= 1'b0;
        end
        else if (stall[0]==`NoStop) begin // shinengxinhao
            ce_reg <= 1'b1;
        end
    end


    assign next_pc = br_e ? br_addr // br_e == 1, next_pc = br_addr 
                   : pc_reg + 32'h4; // br_e == 0, next_pc = pc + 4

    
    assign inst_sram_en = ce_reg; // ID shinengzhiling inst_sram_en = ce_reg
    assign inst_sram_wen = 4'b0; // 
    assign inst_sram_addr = pc_reg; // ID addr = pc_reg
    assign inst_sram_wdata = 32'b0; // 
    assign if_to_id_bus = { //if_to_id_bus zongxian
        ce_reg, //
        pc_reg  //
    };

endmodule